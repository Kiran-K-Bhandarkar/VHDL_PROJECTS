LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FSM_MOORE IS PORT
(
  CLK:    IN STD_LOGIC;
  RST:    IN STD_LOGIC;
  INPUT:  IN STD_LOGIC;
  OUTPUT: OUT STD_LOGIC
);
END ENTITY FSM_MOORE;

ARCHITECTURE BEHAVIORAL OF FSM_MOORE IS
TYPE STATE IS (INIT, A, B, C, D);
SIGNAL CURRENT_STATE, NEXT_STATE: STATE := INIT;
SIGNAL IN_TEMP, OUT_TEMP: STD_LOGIC;

ATTRIBUTE DONT_TOUCH : STRING;
ATTRIBUTE DONT_TOUCH OF  CURRENT_STATE : SIGNAL IS "TRUE";
ATTRIBUTE DONT_TOUCH OF  NEXT_STATE : SIGNAL IS "TRUE";

BEGIN
    IN_TEMP <= INPUT;
	
    -- STATE PROCESS
	PROC_STATE_REG: PROCESS(CLK, RST)
	  BEGIN
		IF RST='1' THEN
		  CURRENT_STATE <= INIT;
		ELSIF RISING_EDGE(CLK) THEN
		  CURRENT_STATE <= NEXT_STATE;
		END IF;
	  END PROCESS PROC_STATE_REG;
	
    --NEXT STATE LOGIC	
	PROC_NSL: PROCESS(CURRENT_STATE, IN_TEMP)
	  BEGIN
		NEXT_STATE <= CURRENT_STATE;
		CASE(CURRENT_STATE) IS
		   WHEN INIT => 
			  IF IN_TEMP = '1' THEN
				NEXT_STATE <= A;
			  END IF;
			  
		   WHEN A => 
			 IF IN_TEMP = '0' THEN
				NEXT_STATE <= B;
			 END IF;
			 
		   WHEN B => 
			 IF IN_TEMP = '1' THEN
				NEXT_STATE <= C;
			ELSE
				NEXT_STATE <= INIT;
			 END IF;
			 
		   WHEN C => 
			 IF IN_TEMP = '0' THEN
				NEXT_STATE <= D;
			 ELSE
				NEXT_STATE <= A;
			 END IF;  
			 
		   WHEN D => 
			 IF IN_TEMP = '1' THEN
				NEXT_STATE <= A;
			 ELSE
			   NEXT_STATE <= INIT;
			 END IF;
		 END CASE;
	END PROCESS PROC_NSL;	 

	-- OUTPUT PROCESS
	PROC_OUT: PROCESS(CURRENT_STATE)
	BEGIN
	  OUT_TEMP <= '0';
	  CASE(CURRENT_STATE) IS
		WHEN D => 
		  OUT_TEMP <= '1';
		WHEN OTHERS =>
		  OUT_TEMP <= '0';
	  END CASE;
	END PROCESS PROC_OUT;
	
	OUTPUT <= OUT_TEMP;
END BEHAVIORAL;
