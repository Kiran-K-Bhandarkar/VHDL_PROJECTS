LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FSM_TB IS 
END ENTITY FSM_TB;

ARCHITECTURE BEHAVIORAL OF FSM_TB IS
SIGNAL CLK, RST, INPUT, OUTPUT: STD_LOGIC;
CONSTANT T: TIME := 5 NS;

BEGIN
  UUT: ENTITY WORK.FSM_MEALY
    PORT MAP
	  (CLK => CLK, RST => RST, INPUT => INPUT, OUTPUT => OUTPUT);
	  
  CLOCK_PROCESS: PROCESS 
    BEGIN
	  CLK <= '0';
	  WAIT FOR T/2;
	  CLK <= '1';
	  WAIT FOR T/2;
	END PROCESS CLOCK_PROCESS;
	
  TEST_PROCESS: PROCESS 
    BEGIN
	  WAIT FOR T;
	  INPUT <= '1';
	  WAIT FOR T;
	  INPUT <= '0';
	  WAIT FOR T;
	  INPUT <= '1';
	  WAIT FOR T;
	  INPUT <= '0';
	  WAIT FOR T;
	  
	  INPUT <= '1';
	  WAIT FOR T;
	  INPUT <= '0';
	  WAIT FOR T;
	  INPUT <= '1';
	  WAIT FOR T;
	  INPUT <= '1';
	  WAIT FOR T;
	   
	  INPUT <= '1';
	  WAIT FOR T;
	  INPUT <= '0';
	  WAIT FOR T;
	  INPUT <= '1';
	  WAIT FOR T;
	  INPUT <= '0';
	  
	  WAIT;
	  END PROCESS TEST_PROCESS;
END BEHAVIORAL;
