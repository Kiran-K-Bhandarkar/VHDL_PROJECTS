LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FSM_MEALY IS PORT 
(
  CLK:    IN STD_LOGIC;
  RST:    IN STD_LOGIC;
  INPUT:  IN STD_LOGIC;
  OUTPUT: OUT STD_LOGIC
);
END ENTITY FSM_MEALY;

ARCHITECTURE BEHAVIORAL OF FSM_MEALY IS 
TYPE STATE IS (INIT, A, B, C);
SIGNAL CURRENT_STATE, NEXT_STATE: STATE := INIT;

SIGNAL OUT_TEMP, IN_TEMP: STD_LOGIC;

BEGIN 
    IN_TEMP <= INPUT;

    -- STATE PROCESS
	PROC_STATE_REG: PROCESS(CLK, RST)
	  BEGIN
	    IF RST='1' THEN
		  CURRENT_STATE <= INIT;
		ELSIF RISING_EDGE(CLK) THEN
          CURRENT_STATE <= NEXT_STATE;
		END IF;
	END PROCESS PROC_STATE_REG;
	
	-- NEXT STATE LOGIC
	PROC_NSL: PROCESS(CURRENT_STATE, IN_TEMP)
	  BEGIN
       OUT_TEMP <= '0';
	   
	   CASE(CURRENT_STATE) IS
	     WHEN INIT =>
		   IF IN_TEMP = '1' THEN
		     NEXT_STATE <= A;
		   END IF;
		 
		 WHEN A => 
		   IF IN_TEMP = '0' THEN
		     NEXT_STATE <= B;
		   END IF;
		 
		 WHEN B =>
		   IF IN_TEMP = '1' THEN 
		     NEXT_STATE <= C;
		   ELSE
		     NEXT_STATE <= INIT;
		   END IF;
		 
		 WHEN C =>
		   IF IN_TEMP = '0' THEN
		     NEXT_STATE <= INIT;
			 OUT_TEMP   <= '1';
		   ELSE
		     NEXT_STATE <= A;
		   END IF;
		END CASE;
	END PROCESS PROC_NSL;
	
	-- OUTPUT PROCESS SYNC WITH CLK
	PROC_OUT: PROCESS(CLK)
	BEGIN
	  IF RISING_EDGE(CLK) THEN
	    OUTPUT <= OUT_TEMP;
	  END IF;
	END PROCESS PROC_OUT;
END BEHAVIORAL;  
	
	
